library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity main_controller is
	generic(
		
	);
	port(
		CLK			:	in std_logic
	);
end entity;

architecture rtl of main_controller is
	
begin

	

end rtl;